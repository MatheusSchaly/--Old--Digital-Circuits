library verilog;
use verilog.vl_types.all;
entity Process_Test_vlg_sample_tst is
    port(
        Clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Process_Test_vlg_sample_tst;
