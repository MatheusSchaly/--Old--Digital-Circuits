library verilog;
use verilog.vl_types.all;
entity FSM_vlg_vec_tst is
end FSM_vlg_vec_tst;
