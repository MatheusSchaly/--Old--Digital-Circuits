library verilog;
use verilog.vl_types.all;
entity Topo_vlg_vec_tst is
end Topo_vlg_vec_tst;
