library verilog;
use verilog.vl_types.all;
entity topo_vlg_check_tst is
    port(
        LEDR            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end topo_vlg_check_tst;
