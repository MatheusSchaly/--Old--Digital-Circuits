library verilog;
use verilog.vl_types.all;
entity top_calc_vlg_vec_tst is
end top_calc_vlg_vec_tst;
