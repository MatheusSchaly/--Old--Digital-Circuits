library verilog;
use verilog.vl_types.all;
entity Process_Test_vlg_check_tst is
    port(
        Result          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Process_Test_vlg_check_tst;
