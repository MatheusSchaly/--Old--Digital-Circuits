library verilog;
use verilog.vl_types.all;
entity topo_vlg_vec_tst is
end topo_vlg_vec_tst;
