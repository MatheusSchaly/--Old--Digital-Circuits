library verilog;
use verilog.vl_types.all;
entity Process_Test_vlg_vec_tst is
end Process_Test_vlg_vec_tst;
