library verilog;
use verilog.vl_types.all;
entity halfadder_vlg_vec_tst is
end halfadder_vlg_vec_tst;
